-----------------------------------------------------
-- Instruction data_mem entity
-- 
-- Contains all the instructions to be run.
-- 
-- data_mem is kept in rows of 32 bits to represent 32-bit
-- registers.
-- 
-- This component initially reads from the file
-- 'instructions.txt' and saves it into a 2d array.
-- 
-- This component takes in a 32-bit address and returns
-- the instruction at that address.
------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity Inst_Mem is
	port (
                CLK         : in STD_LOGIC;
                Load        : in STD_LOGIC;
                last_instr_address  : out STD_LOGIC_VECTOR (31 downto 0);
		Address     : in STD_LOGIC_VECTOR (31 downto 0);
		Instruction : out STD_LOGIC_VECTOR (31 downto 0)
	);
end Inst_Mem;


architecture behavioral of Inst_Mem is	  

    -- 256 byte instruction data_mem (64 rows * 4 bytes/row)
    type mem_array is array(0 to 63) of STD_LOGIC_VECTOR (31 downto 0);
    signal data_mem: mem_array := (
        "00000000000000000000000000000000", -- initialize data data_mem
        "00000000000000000000000000000000", -- mem 1
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000", -- mem 10 
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",  
        "00000000000000000000000000000000", -- mem 20
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000", -- mem 30
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000", -- mem 40
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000", -- mem 50
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000", 
        "00000000000000000000000000000000", -- mem 60
        "00000000000000000000000000000000",
        "00000000000000000000000000000000",
        "00000000000000000000000000000000"
    );

    begin
       MEM_Process: process(CLK)
         begin
            if (Load = '1') then
           --------------------------
--Project1 test
--------------------------
		data_mem(0) <= "00000000000000000100000000100101" ;--00004025
		data_mem(1) <= "10001100000011010000000000110000" ;--8C0D0030
		data_mem(2) <= "10001100000110000000000000110100" ;--8C180034
		data_mem(3) <= "10001100000110010000000000111000" ;--8C190038
		data_mem(4) <= "00000000000110000101000000100000" ;--00185020
		data_mem(5) <= "10101101000010100000000000000000" ;--AD0A0000
		data_mem(6) <= "10101101000010100000000000000100" ;--AD0A0004  -- true
		data_mem(7) <= "00000001101110000100100000100010" ;--01B84822 --true
		data_mem(8) <= "00000001001110000100100000100010" ;--01384822 -- true
		data_mem(9) <= "10001101000010110000000000000000" ;--8D0B0000 -- start loop
		data_mem(10) <= "10001101000011000000000000000100" ;--8D0C0004
		data_mem(11) <= "00000001011011000101000000100000" ;--016C5020--add true
		data_mem(12) <= "10101101000010100000000000001000" ;--AD0A0008-- store memory true
		data_mem(13) <= "00000001000110010100000000100000" ;--01194020 -- increment memory location 
		data_mem(14) <= "00000001001110000100100000100010" ;--01384822 -- decrement loop counter
		data_mem(15) <= "00000000000010010000100000101010" ;--0009082A -- SLT true
		data_mem(16) <= "00010000001000000000000000000001" ;--10200001 --Branch to exit (18)
		data_mem(17) <= "00001000000000000000000000001001" ;--08000009--Jump to 9 
		data_mem(18) <= "00000000000001000010000000100100" ;--00042024-- and
		data_mem(19) <= "00000000000011010010100000100000" ;--000D2820-- add to register 5
		data_mem(20) <= "00001000000000000000000000010110" ;--08000016-- jump to output (22)
		data_mem(21) <= "00000000000110001000000000100010" ;--00188022-- SUB   Final result 1 not -1 because t8 (reg 24) is -1
		data_mem(22) <= "00000001000000000100000000100100" ;--01004024-- register 8=0
		data_mem(23) <= "00000001000010000100100000100000" ;--01084820--  reg 9 = 2* reg8 
		data_mem(24) <= "00000001001010010100100000100000" ;--01294820 -- reg 9 = 2*reg9
		data_mem(25) <= "00000000100010010101000000100000" ;--00895020-- reg 10 = reg9 +reg8
		data_mem(26) <= "10001101010100000000000000000000" ;--8D500000 -- lw reg 16 from memory
		data_mem(27) <= "00000001000110000100000000100000" ;--01184020 -- increment reg 8
		data_mem(28) <= "00000001000001010000100000101010" ;--0105082A -- SLT result into reg 1
		data_mem(29) <= "00010100001000001111111111111001" ;--1420FFF9 -- BNE address for 23
		data_mem(30) <= "00000000000000001100000000100111" ;--0000C027 -- NOR 0,0 set Reg 24 to 1's
		data_mem(31) <= "00000010000110001000000000100111" ;--02188027 -- NOR Reg 16 ,Reg 24 (rest reg16)
		data_mem(32) <= "00001000000000000000000000010101" ;--08000015 -- jump to 21
                last_instr_address <= std_logic_vector(to_unsigned((32)*4, last_instr_address'length));

	end if;

           if(falling_edge(CLK)) then
               --if (Load = '1') then
                  --data_mem(to_integer(unsigned(Address(31 downto 2))))<= Write_Inst;
               --end if;
           end if;
        end process;
 
        -- Since the registers are in multiples of 4 bytes, we can ignore the last two bits
        instruction <= data_mem(to_integer(unsigned(Address(31 downto 2))));

end behavioral;